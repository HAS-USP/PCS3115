module solucao (m, inta, intb, intc, intd, sa, sb, sc, sd, y);
    // Preencha com sua solução aqui

endmodule
// Não inclua os módulos na sua solução!
// O juiz contém os módulos codprisimples e muxsimples fornecidos com este arquivo